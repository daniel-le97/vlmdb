module lmdb

pub type Mdb_filehandle_t = voidptr
