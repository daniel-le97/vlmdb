module vlmdb

pub type Mdb_filehandle_t = voidptr
